module cardinal_cmp #(

)(
    input 
);

//
nic_pe_module npm0(
    .clk(),
    .reset(),
    .net_so(),
    .net_ro(),
    .net_do(),
    .net_polarity(),
    .net_si(),
    .net_ri(),
    .net_di()
);

endmodule